//A program block that creates the environment and initiate the stimulus

program test();
  
  //declare environment handle
  
  initial begin
    //create environment
    
    //initiate the stimulus by calling run of env

  end

endprogram
